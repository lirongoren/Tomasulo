http://code.google.com/p/tomasulo/source/browse/trunk/src/?r=15